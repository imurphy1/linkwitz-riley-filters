*Shelf Filter Testing

.INCLUDE ../Library/Linkwitz-Riley.lib

***Input***
Vin 1 0 ac 1

***Filters***
X1 1 2 0 LR-SLPnon PARAMS: f1 = 300
X2 1 3 0 LR-SLPinv PARAMS: f1 = 300 g2 = 0.707 g1 = 1.414 Switch = 1
X3 1 4 0 LR-SHPnon PARAMS: f2 = 300 g2 = 1.414 Switch = 1
X4 1 5 0 LR-SHPinv PARAMS: f2 = 300 g2 = 1.414 g1 = 0.707 Switch = 1

***Loads***
Rload0 2 0 1meg
Rload1 3 0 1meg
Rload2 4 0 1meg
Rload3 5 0 1meg

.AC dec 100 10 50k
.PROBE V(1) V(2) V(3) V(4) V(5)
.END
