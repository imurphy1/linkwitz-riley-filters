*Buffer Testing

.INCLUDE ../Library/Linkwitz-Riley.lib

***Input***
Vin 1 0 ac 1

***Filters***
X1 1 2 0 LR-NTC1 PARAMS:
X2 1 3 0 LR-NTC2 PARAMS:
X3 1 4 0 LR-NTC3 PARAMS:

***Loads***
Rload0 2 0 1meg
Rload1 3 0 1meg
Rload2 4 0 1meg

.AC dec 100 10 50k
.PROBE V(1) V(2) V(3) V(4)
.END
