*Delay Correction Testing

.INCLUDE ../Library/Linkwitz-Riley.lib

***Input***
Vin 1 0 ac 1

***Filters***
Xd1 1 2 0 LR-D1 PARAMS: f0 = 2500 Switch = 1
Xd2 1 3 0 LR-D2 PARAMS: f0 = 2500 Switch = 1 Ccutoff = 220p

***Loads***
Rload0 2 0 10k
Rload1 3 0 10k

.AC dec 100 10 50000k
.PROBE V(1) V(2) V(3)
.END
